module csa_8 (
  input logic [7:0] a, b,
  input logic cin,
  output logic [7:0] sum,
  output logic cout
);

//do name port association 
logic [3:0] sum1;
logic c0;

adder_4 adder1(.A(a[3:0]), .B(b[3:0]), .cin(cin), .sum(sum1), .cout(c0));


logic [3:0] sum2, sum3;
logic c7_2, c7_3;

//the two parallel adders that compute with both carry 0 and 1
adder_4 adder2(.A(a[7:4]), .B(b[7:4]), .cin(1'b0), .sum(sum2), .cout(c7_2));
adder_4 adder3(.A(a[7:4]), .B(b[7:4]), .cin(1'b1), .sum(sum3), .cout(c7_3));

logic [3:0] s_result;

//first mux for the sum output
always_comb begin 
    s_result = 4'd0;  
    case(c0)
      1'b0: s_result = sum2;
      1'b1: s_result = sum3;
    default: s_result = 4'd0;  
    endcase
end

logic final_carry;

//second mux for the carry 
always_comb begin 
    final_carry = 1'b0;  
    case(c0)
      1'b0: final_carry = c7_2;
      1'b1: final_carry = c7_3;
    default: final_carry = 1'b0;  
    endcase
end

assign cout = final_carry;
assign sum [3:0] = sum1;
assign sum[7:4] = s_result;


endmodule
