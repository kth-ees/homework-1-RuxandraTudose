module csa_8_tb;

  // Inputs
  logic [7:0] a;
  logic [7:0] b;
  logic [7:0] sum;
  logic cin;
  logic cout;

  csa_8 uut (
    .a(a),
    .b(b),
    .sum(sum),
    .cin(cin),
    .cout(cout)
  );

  /* initial begin 
    for(int i = 0; i < 5; i ++) begin
        a = $urandom;
        b = $urandom;
        #10ns;
    end    

  end*/

  initial begin
        a = 8'd33;
        b = 8'd100;
        cin = 1'b0;
  end  
endmodule  

  
  

