module bin2gray (
  input logic [3:0] binary,
  output logic [3:0] gray
);
  // …
  // Add your description here
  // …


  //use 4 MUXES - control singnal Binary values 
  //connect the muxes to the GREY code values 
endmodule
